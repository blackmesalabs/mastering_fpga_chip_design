always @( posedge clk ) begin
  a <= b;
end
