module top
(
  input  wire bd_rx,
  output wire bd_tx
);// module top

  assign bd_tx = bd_rx;
endmodule // top.v
