 reg  foo = 0;
always @ ( posedge clk ) begin
 foo <= bar;
end
