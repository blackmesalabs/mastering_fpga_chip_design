library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
entity rom_font is
port
(
  clk    : in std_logic;
  ck_en  : in std_logic;
  a_addr : in std_logic_vector(11 downto 0);
  a_data : out std_logic_vector(7 downto 0);
  b_addr : in std_logic_vector(11 downto 0);
  b_data : out std_logic_vector(7 downto 0) 
);
end rom_font;
architecture rtl of rom_font is
type rom_type is array (0 to 4095) of std_logic_vector(7 downto 0);
 constant rom : rom_type := (
------ 0
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 1
  "00000000",
  "00000000",
  "01111110",
  "10000001",
  "10100101",
  "10000001",
  "10000001",
  "10111101",
  "10011001",
  "10000001",
  "10000001",
  "01111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 2
  "00000000",
  "00000000",
  "01111110",
  "11111111",
  "11011011",
  "11111111",
  "11111111",
  "11000011",
  "11100111",
  "11111111",
  "11111111",
  "01111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 3
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "01101100",
  "11111110",
  "11111110",
  "11111110",
  "11111110",
  "01111100",
  "00111000",
  "00010000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 4
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00010000",
  "00111000",
  "01111100",
  "11111110",
  "01111100",
  "00111000",
  "00010000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 5
  "00000000",
  "00000000",
  "00000000",
  "00011000",
  "00111100",
  "00111100",
  "11100111",
  "11100111",
  "11100111",
  "00011000",
  "00011000",
  "00111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 6
  "00000000",
  "00000000",
  "00000000",
  "00011000",
  "00111100",
  "01111110",
  "11111111",
  "11111111",
  "01111110",
  "00011000",
  "00011000",
  "00111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 7
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00011000",
  "00111100",
  "00111100",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 8
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11100111",
  "11000011",
  "11000011",
  "11100111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
------ 9
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00111100",
  "01100110",
  "01000010",
  "01000010",
  "01100110",
  "00111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 10
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11000011",
  "10011001",
  "10111101",
  "10111101",
  "10011001",
  "11000011",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
------ 11
  "00000000",
  "00000000",
  "00011110",
  "00001110",
  "00011010",
  "00110010",
  "01111000",
  "11001100",
  "11001100",
  "11001100",
  "11001100",
  "01111000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 12
  "00000000",
  "00000000",
  "00111100",
  "01100110",
  "01100110",
  "01100110",
  "01100110",
  "00111100",
  "00011000",
  "01111110",
  "00011000",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 13
  "00000000",
  "00000000",
  "00111111",
  "00110011",
  "00111111",
  "00110000",
  "00110000",
  "00110000",
  "00110000",
  "01110000",
  "11110000",
  "11100000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 14
  "00000000",
  "00000000",
  "01111111",
  "01100011",
  "01111111",
  "01100011",
  "01100011",
  "01100011",
  "01100011",
  "01100111",
  "11100111",
  "11100110",
  "11000000",
  "00000000",
  "00000000",
  "00000000",
------ 15
  "00000000",
  "00000000",
  "00000000",
  "00011000",
  "00011000",
  "11011011",
  "00111100",
  "11100111",
  "00111100",
  "11011011",
  "00011000",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 16
  "00000000",
  "10000000",
  "11000000",
  "11100000",
  "11110000",
  "11111000",
  "11111110",
  "11111000",
  "11110000",
  "11100000",
  "11000000",
  "10000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 17
  "00000000",
  "00000010",
  "00000110",
  "00001110",
  "00011110",
  "00111110",
  "11111110",
  "00111110",
  "00011110",
  "00001110",
  "00000110",
  "00000010",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 18
  "00000000",
  "00000000",
  "00011000",
  "00111100",
  "01111110",
  "00011000",
  "00011000",
  "00011000",
  "01111110",
  "00111100",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 19
  "00000000",
  "00000000",
  "01100110",
  "01100110",
  "01100110",
  "01100110",
  "01100110",
  "01100110",
  "01100110",
  "00000000",
  "01100110",
  "01100110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 20
  "00000000",
  "00000000",
  "01111111",
  "11011011",
  "11011011",
  "11011011",
  "01111011",
  "00011011",
  "00011011",
  "00011011",
  "00011011",
  "00011011",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 21
  "00000000",
  "01111100",
  "11000110",
  "01100000",
  "00111000",
  "01101100",
  "11000110",
  "11000110",
  "01101100",
  "00111000",
  "00001100",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
------ 22
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11111110",
  "11111110",
  "11111110",
  "11111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 23
  "00000000",
  "00000000",
  "00011000",
  "00111100",
  "01111110",
  "00011000",
  "00011000",
  "00011000",
  "01111110",
  "00111100",
  "00011000",
  "01111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 24
  "00000000",
  "00000000",
  "00011000",
  "00111100",
  "01111110",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 25
  "00000000",
  "00000000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "01111110",
  "00111100",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 26
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00011000",
  "00001100",
  "11111110",
  "00001100",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 27
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00110000",
  "01100000",
  "11111110",
  "01100000",
  "00110000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 28
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11000000",
  "11000000",
  "11000000",
  "11111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 29
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00100100",
  "01100110",
  "11111111",
  "01100110",
  "00100100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 30
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00010000",
  "00111000",
  "00111000",
  "01111100",
  "01111100",
  "11111110",
  "11111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 31
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11111110",
  "11111110",
  "01111100",
  "01111100",
  "00111000",
  "00111000",
  "00010000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 32
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 33
  "00000000",
  "00000000",
  "00011000",
  "00111100",
  "00111100",
  "00111100",
  "00011000",
  "00011000",
  "00011000",
  "00000000",
  "00011000",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 34
  "00000000",
  "01100110",
  "01100110",
  "01100110",
  "00100100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 35
  "00000000",
  "00000000",
  "00000000",
  "01101100",
  "01101100",
  "11111110",
  "01101100",
  "01101100",
  "01101100",
  "11111110",
  "01101100",
  "01101100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 36
  "00011000",
  "00011000",
  "01111100",
  "11000110",
  "11000010",
  "11000000",
  "01111100",
  "00000110",
  "00000110",
  "10000110",
  "11000110",
  "01111100",
  "00011000",
  "00011000",
  "00000000",
  "00000000",
------ 37
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11000010",
  "11000110",
  "00001100",
  "00011000",
  "00110000",
  "01100000",
  "11000110",
  "10000110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 38
  "00000000",
  "00000000",
  "00111000",
  "01101100",
  "01101100",
  "00111000",
  "01110110",
  "11011100",
  "11001100",
  "11001100",
  "11001100",
  "01110110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 39
  "00000000",
  "00110000",
  "00110000",
  "00110000",
  "01100000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 40
  "00000000",
  "00000000",
  "00001100",
  "00011000",
  "00110000",
  "00110000",
  "00110000",
  "00110000",
  "00110000",
  "00110000",
  "00011000",
  "00001100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 41
  "00000000",
  "00000000",
  "00110000",
  "00011000",
  "00001100",
  "00001100",
  "00001100",
  "00001100",
  "00001100",
  "00001100",
  "00011000",
  "00110000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 42
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "01100110",
  "00111100",
  "11111111",
  "00111100",
  "01100110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 43
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00011000",
  "00011000",
  "01111110",
  "00011000",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 44
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00011000",
  "00011000",
  "00011000",
  "00110000",
  "00000000",
  "00000000",
  "00000000",
------ 45
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "01111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 46
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00011000",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 47
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000010",
  "00000110",
  "00001100",
  "00011000",
  "00110000",
  "01100000",
  "11000000",
  "10000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 48
  "00000000",
  "00000000",
  "01111100",
  "11000110",
  "11000110",
  "11001110",
  "11011110",
  "11110110",
  "11100110",
  "11000110",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 49
  "00000000",
  "00000000",
  "00011000",
  "00111000",
  "01111000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "01111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 50
  "00000000",
  "00000000",
  "01111100",
  "11000110",
  "00000110",
  "00001100",
  "00011000",
  "00110000",
  "01100000",
  "11000000",
  "11000110",
  "11111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 51
  "00000000",
  "00000000",
  "01111100",
  "11000110",
  "00000110",
  "00000110",
  "00111100",
  "00000110",
  "00000110",
  "00000110",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 52
  "00000000",
  "00000000",
  "00001100",
  "00011100",
  "00111100",
  "01101100",
  "11001100",
  "11111110",
  "00001100",
  "00001100",
  "00001100",
  "00011110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 53
  "00000000",
  "00000000",
  "11111110",
  "11000000",
  "11000000",
  "11000000",
  "11111100",
  "00000110",
  "00000110",
  "00000110",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 54
  "00000000",
  "00000000",
  "00111000",
  "01100000",
  "11000000",
  "11000000",
  "11111100",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 55
  "00000000",
  "00000000",
  "11111110",
  "11000110",
  "00000110",
  "00000110",
  "00001100",
  "00011000",
  "00110000",
  "00110000",
  "00110000",
  "00110000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 56
  "00000000",
  "00000000",
  "01111100",
  "11000110",
  "11000110",
  "11000110",
  "01111100",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 57
  "00000000",
  "00000000",
  "01111100",
  "11000110",
  "11000110",
  "11000110",
  "01111110",
  "00000110",
  "00000110",
  "00000110",
  "00001100",
  "01111000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 58
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00011000",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00011000",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 59
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00011000",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00011000",
  "00011000",
  "00110000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 60
  "00000000",
  "00000000",
  "00000000",
  "00000110",
  "00001100",
  "00011000",
  "00110000",
  "01100000",
  "00110000",
  "00011000",
  "00001100",
  "00000110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 61
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "01111110",
  "00000000",
  "00000000",
  "01111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 62
  "00000000",
  "00000000",
  "00000000",
  "01100000",
  "00110000",
  "00011000",
  "00001100",
  "00000110",
  "00001100",
  "00011000",
  "00110000",
  "01100000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 63
  "00000000",
  "00000000",
  "01111100",
  "11000110",
  "11000110",
  "00001100",
  "00011000",
  "00011000",
  "00011000",
  "00000000",
  "00011000",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 64
  "00000000",
  "00000000",
  "01111100",
  "11000110",
  "11000110",
  "11000110",
  "11011110",
  "11011110",
  "11011110",
  "11011100",
  "11000000",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 65
  "00000000",
  "00000000",
  "00010000",
  "00111000",
  "01101100",
  "11000110",
  "11000110",
  "11111110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 66
  "00000000",
  "00000000",
  "11111100",
  "01100110",
  "01100110",
  "01100110",
  "01111100",
  "01100110",
  "01100110",
  "01100110",
  "01100110",
  "11111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 67
  "00000000",
  "00000000",
  "00111100",
  "01100110",
  "11000010",
  "11000000",
  "11000000",
  "11000000",
  "11000000",
  "11000010",
  "01100110",
  "00111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 68
  "00000000",
  "00000000",
  "11111000",
  "01101100",
  "01100110",
  "01100110",
  "01100110",
  "01100110",
  "01100110",
  "01100110",
  "01101100",
  "11111000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 69
  "00000000",
  "00000000",
  "11111110",
  "01100110",
  "01100010",
  "01101000",
  "01111000",
  "01101000",
  "01100000",
  "01100010",
  "01100110",
  "11111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 70
  "00000000",
  "00000000",
  "11111110",
  "01100110",
  "01100010",
  "01101000",
  "01111000",
  "01101000",
  "01100000",
  "01100000",
  "01100000",
  "11110000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 71
  "00000000",
  "00000000",
  "00111100",
  "01100110",
  "11000010",
  "11000000",
  "11000000",
  "11011110",
  "11000110",
  "11000110",
  "01100110",
  "00111010",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 72
  "00000000",
  "00000000",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11111110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 73
  "00000000",
  "00000000",
  "00111100",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 74
  "00000000",
  "00000000",
  "00011110",
  "00001100",
  "00001100",
  "00001100",
  "00001100",
  "00001100",
  "11001100",
  "11001100",
  "11001100",
  "01111000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 75
  "00000000",
  "00000000",
  "11100110",
  "01100110",
  "01100110",
  "01101100",
  "01111000",
  "01111000",
  "01101100",
  "01100110",
  "01100110",
  "11100110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 76
  "00000000",
  "00000000",
  "11110000",
  "01100000",
  "01100000",
  "01100000",
  "01100000",
  "01100000",
  "01100000",
  "01100010",
  "01100110",
  "11111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 77
  "00000000",
  "00000000",
  "11000011",
  "11100111",
  "11111111",
  "11111111",
  "11011011",
  "11000011",
  "11000011",
  "11000011",
  "11000011",
  "11000011",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 78
  "00000000",
  "00000000",
  "11000110",
  "11100110",
  "11110110",
  "11111110",
  "11011110",
  "11001110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 79
  "00000000",
  "00000000",
  "01111100",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 80
  "00000000",
  "00000000",
  "11111100",
  "01100110",
  "01100110",
  "01100110",
  "01111100",
  "01100000",
  "01100000",
  "01100000",
  "01100000",
  "11110000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 81
  "00000000",
  "00000000",
  "01111100",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11010110",
  "11011110",
  "01111100",
  "00001100",
  "00001110",
  "00000000",
  "00000000",
------ 82
  "00000000",
  "00000000",
  "11111100",
  "01100110",
  "01100110",
  "01100110",
  "01111100",
  "01101100",
  "01100110",
  "01100110",
  "01100110",
  "11100110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 83
  "00000000",
  "00000000",
  "01111100",
  "11000110",
  "11000110",
  "01100000",
  "00111000",
  "00001100",
  "00000110",
  "11000110",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 84
  "00000000",
  "00000000",
  "11111111",
  "11011011",
  "10011001",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 85
  "00000000",
  "00000000",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 86
  "00000000",
  "00000000",
  "11000011",
  "11000011",
  "11000011",
  "11000011",
  "11000011",
  "11000011",
  "11000011",
  "01100110",
  "00111100",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 87
  "00000000",
  "00000000",
  "11000011",
  "11000011",
  "11000011",
  "11000011",
  "11000011",
  "11011011",
  "11011011",
  "11111111",
  "01100110",
  "01100110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 88
  "00000000",
  "00000000",
  "11000011",
  "11000011",
  "01100110",
  "00111100",
  "00011000",
  "00011000",
  "00111100",
  "01100110",
  "11000011",
  "11000011",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 89
  "00000000",
  "00000000",
  "11000011",
  "11000011",
  "11000011",
  "01100110",
  "00111100",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 90
  "00000000",
  "00000000",
  "11111111",
  "11000011",
  "10000110",
  "00001100",
  "00011000",
  "00110000",
  "01100000",
  "11000001",
  "11000011",
  "11111111",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 91
  "00000000",
  "00000000",
  "00111100",
  "00110000",
  "00110000",
  "00110000",
  "00110000",
  "00110000",
  "00110000",
  "00110000",
  "00110000",
  "00111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 92
  "00000000",
  "00000000",
  "00000000",
  "10000000",
  "11000000",
  "11100000",
  "01110000",
  "00111000",
  "00011100",
  "00001110",
  "00000110",
  "00000010",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 93
  "00000000",
  "00000000",
  "00111100",
  "00001100",
  "00001100",
  "00001100",
  "00001100",
  "00001100",
  "00001100",
  "00001100",
  "00001100",
  "00111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 94
  "00010000",
  "00111000",
  "01101100",
  "11000110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 95
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11111111",
  "00000000",
  "00000000",
------ 96
  "00110000",
  "00110000",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 97
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "01111000",
  "00001100",
  "01111100",
  "11001100",
  "11001100",
  "11001100",
  "01110110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 98
  "00000000",
  "00000000",
  "11100000",
  "01100000",
  "01100000",
  "01111000",
  "01101100",
  "01100110",
  "01100110",
  "01100110",
  "01100110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 99
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "01111100",
  "11000110",
  "11000000",
  "11000000",
  "11000000",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 100
  "00000000",
  "00000000",
  "00011100",
  "00001100",
  "00001100",
  "00111100",
  "01101100",
  "11001100",
  "11001100",
  "11001100",
  "11001100",
  "01110110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 101
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "01111100",
  "11000110",
  "11111110",
  "11000000",
  "11000000",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 102
  "00000000",
  "00000000",
  "00111000",
  "01101100",
  "01100100",
  "01100000",
  "11110000",
  "01100000",
  "01100000",
  "01100000",
  "01100000",
  "11110000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 103
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "01110110",
  "11001100",
  "11001100",
  "11001100",
  "11001100",
  "11001100",
  "01111100",
  "00001100",
  "11001100",
  "01111000",
  "00000000",
------ 104
  "00000000",
  "00000000",
  "11100000",
  "01100000",
  "01100000",
  "01101100",
  "01110110",
  "01100110",
  "01100110",
  "01100110",
  "01100110",
  "11100110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 105
  "00000000",
  "00000000",
  "00011000",
  "00011000",
  "00000000",
  "00111000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 106
  "00000000",
  "00000000",
  "00000110",
  "00000110",
  "00000000",
  "00001110",
  "00000110",
  "00000110",
  "00000110",
  "00000110",
  "00000110",
  "00000110",
  "01100110",
  "01100110",
  "00111100",
  "00000000",
------ 107
  "00000000",
  "00000000",
  "11100000",
  "01100000",
  "01100000",
  "01100110",
  "01101100",
  "01111000",
  "01111000",
  "01101100",
  "01100110",
  "11100110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 108
  "00000000",
  "00000000",
  "00111000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 109
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11100110",
  "11111111",
  "11011011",
  "11011011",
  "11011011",
  "11011011",
  "11011011",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 110
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11011100",
  "01100110",
  "01100110",
  "01100110",
  "01100110",
  "01100110",
  "01100110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 111
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "01111100",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 112
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11011100",
  "01100110",
  "01100110",
  "01100110",
  "01100110",
  "01100110",
  "01111100",
  "01100000",
  "01100000",
  "11110000",
  "00000000",
------ 113
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "01110110",
  "11001100",
  "11001100",
  "11001100",
  "11001100",
  "11001100",
  "01111100",
  "00001100",
  "00001100",
  "00011110",
  "00000000",
------ 114
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11011100",
  "01110110",
  "01100110",
  "01100000",
  "01100000",
  "01100000",
  "11110000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 115
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "01111100",
  "11000110",
  "01100000",
  "00111000",
  "00001100",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 116
  "00000000",
  "00000000",
  "00010000",
  "00110000",
  "00110000",
  "11111100",
  "00110000",
  "00110000",
  "00110000",
  "00110000",
  "00110110",
  "00011100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 117
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11001100",
  "11001100",
  "11001100",
  "11001100",
  "11001100",
  "11001100",
  "01110110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 118
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11000011",
  "11000011",
  "11000011",
  "11000011",
  "01100110",
  "00111100",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 119
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11000011",
  "11000011",
  "11000011",
  "11011011",
  "11011011",
  "11111111",
  "01100110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 120
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11000011",
  "01100110",
  "00111100",
  "00011000",
  "00111100",
  "01100110",
  "11000011",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 121
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "01111110",
  "00000110",
  "00001100",
  "11111000",
  "00000000",
------ 122
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11111110",
  "11001100",
  "00011000",
  "00110000",
  "01100000",
  "11000110",
  "11111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 123
  "00000000",
  "00000000",
  "00001110",
  "00011000",
  "00011000",
  "00011000",
  "01110000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00001110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 124
  "00000000",
  "00000000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00000000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 125
  "00000000",
  "00000000",
  "01110000",
  "00011000",
  "00011000",
  "00011000",
  "00001110",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "01110000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 126
  "00000000",
  "00000000",
  "01110110",
  "11011100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 127
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00010000",
  "00111000",
  "01101100",
  "11000110",
  "11000110",
  "11000110",
  "11111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 128
  "00000000",
  "00000000",
  "00111100",
  "01100110",
  "11000010",
  "11000000",
  "11000000",
  "11000000",
  "11000010",
  "01100110",
  "00111100",
  "00001100",
  "00000110",
  "01111100",
  "00000000",
  "00000000",
------ 129
  "00000000",
  "00000000",
  "11001100",
  "00000000",
  "00000000",
  "11001100",
  "11001100",
  "11001100",
  "11001100",
  "11001100",
  "11001100",
  "01110110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 130
  "00000000",
  "00001100",
  "00011000",
  "00110000",
  "00000000",
  "01111100",
  "11000110",
  "11111110",
  "11000000",
  "11000000",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 131
  "00000000",
  "00010000",
  "00111000",
  "01101100",
  "00000000",
  "01111000",
  "00001100",
  "01111100",
  "11001100",
  "11001100",
  "11001100",
  "01110110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 132
  "00000000",
  "00000000",
  "11001100",
  "00000000",
  "00000000",
  "01111000",
  "00001100",
  "01111100",
  "11001100",
  "11001100",
  "11001100",
  "01110110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 133
  "00000000",
  "01100000",
  "00110000",
  "00011000",
  "00000000",
  "01111000",
  "00001100",
  "01111100",
  "11001100",
  "11001100",
  "11001100",
  "01110110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 134
  "00000000",
  "00111000",
  "01101100",
  "00111000",
  "00000000",
  "01111000",
  "00001100",
  "01111100",
  "11001100",
  "11001100",
  "11001100",
  "01110110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 135
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00111100",
  "01100110",
  "01100000",
  "01100000",
  "01100110",
  "00111100",
  "00001100",
  "00000110",
  "00111100",
  "00000000",
  "00000000",
  "00000000",
------ 136
  "00000000",
  "00010000",
  "00111000",
  "01101100",
  "00000000",
  "01111100",
  "11000110",
  "11111110",
  "11000000",
  "11000000",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 137
  "00000000",
  "00000000",
  "11000110",
  "00000000",
  "00000000",
  "01111100",
  "11000110",
  "11111110",
  "11000000",
  "11000000",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 138
  "00000000",
  "01100000",
  "00110000",
  "00011000",
  "00000000",
  "01111100",
  "11000110",
  "11111110",
  "11000000",
  "11000000",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 139
  "00000000",
  "00000000",
  "01100110",
  "00000000",
  "00000000",
  "00111000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 140
  "00000000",
  "00011000",
  "00111100",
  "01100110",
  "00000000",
  "00111000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 141
  "00000000",
  "01100000",
  "00110000",
  "00011000",
  "00000000",
  "00111000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 142
  "00000000",
  "11000110",
  "00000000",
  "00010000",
  "00111000",
  "01101100",
  "11000110",
  "11000110",
  "11111110",
  "11000110",
  "11000110",
  "11000110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 143
  "00111000",
  "01101100",
  "00111000",
  "00000000",
  "00111000",
  "01101100",
  "11000110",
  "11000110",
  "11111110",
  "11000110",
  "11000110",
  "11000110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 144
  "00011000",
  "00110000",
  "01100000",
  "00000000",
  "11111110",
  "01100110",
  "01100000",
  "01111100",
  "01100000",
  "01100000",
  "01100110",
  "11111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 145
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "01101110",
  "00111011",
  "00011011",
  "01111110",
  "11011000",
  "11011100",
  "01110111",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 146
  "00000000",
  "00000000",
  "00111110",
  "01101100",
  "11001100",
  "11001100",
  "11111110",
  "11001100",
  "11001100",
  "11001100",
  "11001100",
  "11001110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 147
  "00000000",
  "00010000",
  "00111000",
  "01101100",
  "00000000",
  "01111100",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 148
  "00000000",
  "00000000",
  "11000110",
  "00000000",
  "00000000",
  "01111100",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 149
  "00000000",
  "01100000",
  "00110000",
  "00011000",
  "00000000",
  "01111100",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 150
  "00000000",
  "00110000",
  "01111000",
  "11001100",
  "00000000",
  "11001100",
  "11001100",
  "11001100",
  "11001100",
  "11001100",
  "11001100",
  "01110110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 151
  "00000000",
  "01100000",
  "00110000",
  "00011000",
  "00000000",
  "11001100",
  "11001100",
  "11001100",
  "11001100",
  "11001100",
  "11001100",
  "01110110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 152
  "00000000",
  "00000000",
  "11000110",
  "00000000",
  "00000000",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "01111110",
  "00000110",
  "00001100",
  "01111000",
  "00000000",
------ 153
  "00000000",
  "11000110",
  "00000000",
  "01111100",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 154
  "00000000",
  "11000110",
  "00000000",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 155
  "00000000",
  "00011000",
  "00011000",
  "01111110",
  "11000011",
  "11000000",
  "11000000",
  "11000000",
  "11000011",
  "01111110",
  "00011000",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 156
  "00000000",
  "00111000",
  "01101100",
  "01100100",
  "01100000",
  "11110000",
  "01100000",
  "01100000",
  "01100000",
  "01100000",
  "11100110",
  "11111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 157
  "00000000",
  "00000000",
  "11000011",
  "01100110",
  "00111100",
  "00011000",
  "11111111",
  "00011000",
  "11111111",
  "00011000",
  "00011000",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 158
  "00000000",
  "11111100",
  "01100110",
  "01100110",
  "01111100",
  "01100010",
  "01100110",
  "01101111",
  "01100110",
  "01100110",
  "01100110",
  "11110011",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 159
  "00000000",
  "00001110",
  "00011011",
  "00011000",
  "00011000",
  "00011000",
  "01111110",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "11011000",
  "01110000",
  "00000000",
  "00000000",
------ 160
  "00000000",
  "00011000",
  "00110000",
  "01100000",
  "00000000",
  "01111000",
  "00001100",
  "01111100",
  "11001100",
  "11001100",
  "11001100",
  "01110110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 161
  "00000000",
  "00001100",
  "00011000",
  "00110000",
  "00000000",
  "00111000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 162
  "00000000",
  "00011000",
  "00110000",
  "01100000",
  "00000000",
  "01111100",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 163
  "00000000",
  "00011000",
  "00110000",
  "01100000",
  "00000000",
  "11001100",
  "11001100",
  "11001100",
  "11001100",
  "11001100",
  "11001100",
  "01110110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 164
  "00000000",
  "00000000",
  "01110110",
  "11011100",
  "00000000",
  "11011100",
  "01100110",
  "01100110",
  "01100110",
  "01100110",
  "01100110",
  "01100110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 165
  "01110110",
  "11011100",
  "00000000",
  "11000110",
  "11100110",
  "11110110",
  "11111110",
  "11011110",
  "11001110",
  "11000110",
  "11000110",
  "11000110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 166
  "00000000",
  "00111100",
  "01101100",
  "01101100",
  "00111110",
  "00000000",
  "01111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 167
  "00000000",
  "00111000",
  "01101100",
  "01101100",
  "00111000",
  "00000000",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 168
  "00000000",
  "00000000",
  "00110000",
  "00110000",
  "00000000",
  "00110000",
  "00110000",
  "01100000",
  "11000000",
  "11000110",
  "11000110",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 169
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11111110",
  "11000000",
  "11000000",
  "11000000",
  "11000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 170
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11111110",
  "00000110",
  "00000110",
  "00000110",
  "00000110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 171
  "00000000",
  "11000000",
  "11000000",
  "11000010",
  "11000110",
  "11001100",
  "00011000",
  "00110000",
  "01100000",
  "11001110",
  "10011011",
  "00000110",
  "00001100",
  "00011111",
  "00000000",
  "00000000",
------ 172
  "00000000",
  "11000000",
  "11000000",
  "11000010",
  "11000110",
  "11001100",
  "00011000",
  "00110000",
  "01100110",
  "11001110",
  "10010110",
  "00111110",
  "00000110",
  "00000110",
  "00000000",
  "00000000",
------ 173
  "00000000",
  "00000000",
  "00011000",
  "00011000",
  "00000000",
  "00011000",
  "00011000",
  "00011000",
  "00111100",
  "00111100",
  "00111100",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 174
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00110110",
  "01101100",
  "11011000",
  "01101100",
  "00110110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 175
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11011000",
  "01101100",
  "00110110",
  "01101100",
  "11011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 176
  "00010001",
  "01000100",
  "00010001",
  "01000100",
  "00010001",
  "01000100",
  "00010001",
  "01000100",
  "00010001",
  "01000100",
  "00010001",
  "01000100",
  "00010001",
  "01000100",
  "00010001",
  "01000100",
------ 177
  "01010101",
  "10101010",
  "01010101",
  "10101010",
  "01010101",
  "10101010",
  "01010101",
  "10101010",
  "01010101",
  "10101010",
  "01010101",
  "10101010",
  "01010101",
  "10101010",
  "01010101",
  "10101010",
------ 178
  "11011101",
  "01110111",
  "11011101",
  "01110111",
  "11011101",
  "01110111",
  "11011101",
  "01110111",
  "11011101",
  "01110111",
  "11011101",
  "01110111",
  "11011101",
  "01110111",
  "11011101",
  "01110111",
------ 179
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
------ 180
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "11111000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
------ 181
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "11111000",
  "00011000",
  "11111000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
------ 182
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "11110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
------ 183
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11111110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
------ 184
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11111000",
  "00011000",
  "11111000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
------ 185
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "11110110",
  "00000110",
  "11110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
------ 186
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
------ 187
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11111110",
  "00000110",
  "11110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
------ 188
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "11110110",
  "00000110",
  "11111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 189
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "11111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 190
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "11111000",
  "00011000",
  "11111000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 191
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11111000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
------ 192
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011111",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 193
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "11111111",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 194
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11111111",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
------ 195
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011111",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
------ 196
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11111111",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 197
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "11111111",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
------ 198
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011111",
  "00011000",
  "00011111",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
------ 199
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110111",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
------ 200
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110111",
  "00110000",
  "00111111",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 201
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00111111",
  "00110000",
  "00110111",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
------ 202
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "11110111",
  "00000000",
  "11111111",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 203
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11111111",
  "00000000",
  "11110111",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
------ 204
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110111",
  "00110000",
  "00110111",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
------ 205
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11111111",
  "00000000",
  "11111111",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 206
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "11110111",
  "00000000",
  "11110111",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
------ 207
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "11111111",
  "00000000",
  "11111111",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 208
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "11111111",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 209
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11111111",
  "00000000",
  "11111111",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
------ 210
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11111111",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
------ 211
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00111111",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 212
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011111",
  "00011000",
  "00011111",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 213
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00011111",
  "00011000",
  "00011111",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
------ 214
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00111111",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
------ 215
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "11111111",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
  "00110110",
------ 216
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "11111111",
  "00011000",
  "11111111",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
------ 217
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "11111000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 218
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00011111",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
------ 219
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
------ 220
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
------ 221
  "11110000",
  "11110000",
  "11110000",
  "11110000",
  "11110000",
  "11110000",
  "11110000",
  "11110000",
  "11110000",
  "11110000",
  "11110000",
  "11110000",
  "11110000",
  "11110000",
  "11110000",
  "11110000",
------ 222
  "00001111",
  "00001111",
  "00001111",
  "00001111",
  "00001111",
  "00001111",
  "00001111",
  "00001111",
  "00001111",
  "00001111",
  "00001111",
  "00001111",
  "00001111",
  "00001111",
  "00001111",
  "00001111",
------ 223
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "11111111",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 224
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "01110110",
  "11011100",
  "11011000",
  "11011000",
  "11011000",
  "11011100",
  "01110110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 225
  "00000000",
  "00000000",
  "01111000",
  "11001100",
  "11001100",
  "11001100",
  "11011000",
  "11001100",
  "11000110",
  "11000110",
  "11000110",
  "11001100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 226
  "00000000",
  "00000000",
  "11111110",
  "11000110",
  "11000110",
  "11000000",
  "11000000",
  "11000000",
  "11000000",
  "11000000",
  "11000000",
  "11000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 227
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11111110",
  "01101100",
  "01101100",
  "01101100",
  "01101100",
  "01101100",
  "01101100",
  "01101100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 228
  "00000000",
  "00000000",
  "00000000",
  "11111110",
  "11000110",
  "01100000",
  "00110000",
  "00011000",
  "00110000",
  "01100000",
  "11000110",
  "11111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 229
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "01111110",
  "11011000",
  "11011000",
  "11011000",
  "11011000",
  "11011000",
  "01110000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 230
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "01100110",
  "01100110",
  "01100110",
  "01100110",
  "01100110",
  "01111100",
  "01100000",
  "01100000",
  "11000000",
  "00000000",
  "00000000",
  "00000000",
------ 231
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "01110110",
  "11011100",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 232
  "00000000",
  "00000000",
  "00000000",
  "01111110",
  "00011000",
  "00111100",
  "01100110",
  "01100110",
  "01100110",
  "00111100",
  "00011000",
  "01111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 233
  "00000000",
  "00000000",
  "00000000",
  "00111000",
  "01101100",
  "11000110",
  "11000110",
  "11111110",
  "11000110",
  "11000110",
  "01101100",
  "00111000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 234
  "00000000",
  "00000000",
  "00111000",
  "01101100",
  "11000110",
  "11000110",
  "11000110",
  "01101100",
  "01101100",
  "01101100",
  "01101100",
  "11101110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 235
  "00000000",
  "00000000",
  "00011110",
  "00110000",
  "00011000",
  "00001100",
  "00111110",
  "01100110",
  "01100110",
  "01100110",
  "01100110",
  "00111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 236
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "01111110",
  "11011011",
  "11011011",
  "11011011",
  "01111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 237
  "00000000",
  "00000000",
  "00000000",
  "00000011",
  "00000110",
  "01111110",
  "11011011",
  "11011011",
  "11110011",
  "01111110",
  "01100000",
  "11000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 238
  "00000000",
  "00000000",
  "00011100",
  "00110000",
  "01100000",
  "01100000",
  "01111100",
  "01100000",
  "01100000",
  "01100000",
  "00110000",
  "00011100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 239
  "00000000",
  "00000000",
  "00000000",
  "01111100",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "11000110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 240
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "11111110",
  "00000000",
  "00000000",
  "11111110",
  "00000000",
  "00000000",
  "11111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 241
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00011000",
  "00011000",
  "01111110",
  "00011000",
  "00011000",
  "00000000",
  "00000000",
  "11111111",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 242
  "00000000",
  "00000000",
  "00000000",
  "00110000",
  "00011000",
  "00001100",
  "00000110",
  "00001100",
  "00011000",
  "00110000",
  "00000000",
  "01111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 243
  "00000000",
  "00000000",
  "00000000",
  "00001100",
  "00011000",
  "00110000",
  "01100000",
  "00110000",
  "00011000",
  "00001100",
  "00000000",
  "01111110",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 244
  "00000000",
  "00000000",
  "00001110",
  "00011011",
  "00011011",
  "00011011",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
------ 245
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "00011000",
  "11011000",
  "11011000",
  "11011000",
  "01110000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 246
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00011000",
  "00011000",
  "00000000",
  "01111110",
  "00000000",
  "00011000",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 247
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "01110110",
  "11011100",
  "00000000",
  "01110110",
  "11011100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 248
  "00000000",
  "00111000",
  "01101100",
  "01101100",
  "00111000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 249
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00011000",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 250
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00011000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 251
  "00000000",
  "00001111",
  "00001100",
  "00001100",
  "00001100",
  "00001100",
  "00001100",
  "11101100",
  "01101100",
  "01101100",
  "00111100",
  "00011100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 252
  "00000000",
  "11011000",
  "01101100",
  "01101100",
  "01101100",
  "01101100",
  "01101100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 253
  "00000000",
  "01110000",
  "11011000",
  "00110000",
  "01100000",
  "11001000",
  "11111000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 254
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "01111100",
  "01111100",
  "01111100",
  "01111100",
  "01111100",
  "01111100",
  "01111100",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
------ 255
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000",
  "00000000"
 );

begin

flop_proc : process ( clk )
begin
 if ( clk'event and clk = '1' ) then
   if ( ck_en = '1' ) then
     a_data <= rom( conv_integer( a_addr ) );
     b_data <= rom( conv_integer( b_addr ) );
   end if;
 end if;
end process flop_proc;

end rtl;
